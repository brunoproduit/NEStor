

 
 
 




window new WaveWindow  -name  "Waves for BMG Example Design"
waveform  using  "Waves for BMG Example Design"

      waveform add -signals /end_game_screen1_ram_tb/status
      waveform add -signals /end_game_screen1_ram_tb/end_game_screen1_ram_synth_inst/bmg_port/CLKA
      waveform add -signals /end_game_screen1_ram_tb/end_game_screen1_ram_synth_inst/bmg_port/ADDRA
      waveform add -signals /end_game_screen1_ram_tb/end_game_screen1_ram_synth_inst/bmg_port/DOUTA

console submit -using simulator -wait no "run"
